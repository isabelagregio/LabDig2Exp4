module exp5_fd #(
    parameter TIME = 100_000_000
) (
    input clock,
    input reset,
    input medir,
    input echo,
    input partida_serial,
    input zera_timeout_echo,
    input zera_contador_ascii,
    input reset_circuito,
    input conta_ascii,
    input conta_angulo,
    input conta_timeout_echo,
    output fim_serial,
    output trigger,
    output saida_serial,
    output pronto_medida,
    output pronto_transmissao,
    output [11:0] medida,
    output pwm,
    output timeout_echo,
    output [2:0] db_posicao,
    output db_pwm,
    output [3:0] db_estado_medida,
    output [3:0] db_estado_serial,
    output db_partida_serial,
    output db_conta_ascii,
    output db_conta_timeout_echo,
    output db_conta_angulo,
    output db_pronto_medida,
    output db_pronto_transmissao,
	output dois_segundos
);

    wire [6:0] dados_ascii;
    wire [11:0] s_medida;
    wire [23:0] saida_rom;
    wire [2:0] seletor;
    wire [2:0] posicao_angulo;
    
	assign medida = s_medida;

    tx_serial_7E1 tx_serial (
       .clock(clock),
       .reset(reset),
       .partida(partida_serial), 
       .dados_ascii(dados_ascii),
       .saida_serial(saida_serial), 
       .pronto(pronto_transmissao),
       .db_clock(), 
       .db_tick(),
       .db_partida(),
       .db_saida_serial(),
       .db_estado(db_estado_serial)   
    );

    interface_hcsr04 hcsr04(
        .clock(clock),
        .reset(reset),
        .medir(medir),
        .echo(echo),
        .trigger(trigger),
        .medida(s_medida),
        .pronto(pronto_medida),
        .db_estado(db_estado_medida)
    );

    controle_servo_8 controle_servo (
        .clock(clock),
        .reset(reset),
        .posicao(posicao_angulo),
        .controle(pwm), // pwm ligado no servomotor
        .db_controle(db_pwm), // pwm gerado pra depuração
        .db_posicao(db_posicao)
    );

     mux_8x1_n #(
        .BITS(7)
    ) mux_inst (
        .D7(7'h23),
        .D6({3'b000, s_medida[3:0]} + 7'h30),  
        .D5({3'b000, s_medida[7:4]} + 7'h30),   
        .D4({3'b000, s_medida[11:8]} + 7'h30),
        .D3(7'h2C),
        .D2(saida_rom[6:0]),  // descarte do bit mais significativo
        .D1(saida_rom[14:8]),
        .D0(saida_rom[22:16]),
        .SEL(seletor),
        .MUX_OUT(dados_ascii)
    );

    rom_angulos_8x24 rom (
        .endereco(posicao_angulo), 
        .saida(saida_rom)
    );
  
    contador_m #(  // contador blocos ascii
        .M (8), 
        .N (3)
    ) contador_ascii (
        .clock   (clock     ),
        .zera_as (1'b0      ),
        .zera_s  (zera_contador_ascii ),
        .conta   (conta_ascii),
        .Q       (seletor), 
        .fim     (fim_serial),  
        .meio    (      )
    );

    contador_m #(  // contador angulos
        .M (8), 
        .N (3)
    ) contador_angulos (
        .clock   (clock     ),
        .zera_as (1'b0      ),
        .zera_s  (reset_circuito ),
        .conta   (conta_angulo),
        .Q       (posicao_angulo), 
        .fim     (),  
        .meio    (      )
    );

	   
    contador_m #(   // timer de 2 segundos
        .M (TIME), 
        .N (27)
    ) contador_segundo (
        .clock   (clock     ),
        .zera_as (1'b0      ),
        .zera_s  (reset_circuito ),
        .conta   (1'b1),
        .Q       (), 
        .fim     (dois_segundos),  
        .meio    (      )
    );

    contador_m #(   // timer de 200 milisegundos
        .M (10_000_000), 
        .N (24)
    ) contador_timeout_echo (
        .clock   (clock     ),
        .zera_as (1'b0      ),
        .zera_s  (zera_timeout_echo ),
        .conta   (conta_timeout_echo),
        .Q       (), 
        .fim     (timeout_echo),  
        .meio    (      )
    );
	 
	 
endmodule